module configuration_manager